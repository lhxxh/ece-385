module testbench();

timeunit 10ns;

timeprecision 1ns;

	logic CLK;
	logic RESET;
	logic AES_START;
	logic AES_DONE;
	logic [127:0] AES_KEY;
	logic [127:0] AES_MSG_ENC;
	logic [127:0] AES_MSG_DEC;

always begin : CLOCK_GENERATION
 
 #1 CLK = ~CLK;
 
 end
 
initial begin : CLOCK_INITIALIZATION
	
    CLK = 0;
	
 end
 
 AES tp(.*);
 
 initial begin : TEST_VECTORS
 

 
  RESET = 1;
 
 #2 RESET = 0;
 
 AES_KEY = 128'b00000000000000010000001000000011000001000000010100000110000001110000100000001001000010100000101100001100000011010000111000001111;
 AES_MSG_ENC = 128'b11011010111011000011000001010101110111110000010110001110000111000011100111101000000101001110101001110110111101100111010001111110;
 
 #10 AES_START = 1;
 
 
 
 end

endmodule